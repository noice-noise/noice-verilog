module verilog_tb();
    reg